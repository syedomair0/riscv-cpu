module alu(
	
);

endmodule

module prefix_adder(
	input[15:0] a,
	input[15:0] b
);

// generate signal is a & b
// propogate signal is a | b



endmodule
